library IEEE; 
use IEEE.STD_LOGIC_1164.all;

entity aludec is -- ALU control decoder
  port(funct:      in  STD_LOGIC_VECTOR(5 downto 0);
       aluop:      in  STD_LOGIC_VECTOR(2 downto 0);
       alucontrol: out STD_LOGIC_VECTOR(2 downto 0));
end;

-------------------------------------------------------------------------
-- Elizabeth Roberts, Benjamin Greenwood, Christopher Oriolt and Shane Snediker
-- CS 401 MIPS 4
--Last updated: 3-24-21
-------------------------------------------------------------------------
architecture behave of aludec is
begin
  process(aluop, funct) begin
    case aluop is
      when "000" => alucontrol <= "010"; -- add (for lb/sb/addi)
      when "001" => alucontrol <= "110"; -- sub (for beq)
      when "100" => alucontrol <= "011"; -- SLTi 
      when "101" => alucontrol <= "101"; -- ORI
      when others => case funct is         -- R-type instructions
          when "100000" => alucontrol <= "010"; -- add (for add)
          when "100010" => alucontrol <= "110"; -- subtract (for sub)
          when "100100" => alucontrol <= "000"; -- logical and (for and)
          when "100101" => alucontrol <= "001"; -- logical or (for or)
          when "000000" => alucontrol <= "100"; -- shift left logical
          when "000010" => alucontrol <= "111"; -- shift right logical
          when others   => alucontrol <= "---"; -- should never happen
        end case;
    end case;
  end process;
end;

